`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "memory.v"
`include "mem_assertion.sv"
`include "mem_intf.sv"
`include "mem_tx.sv"
`include "mem_cov.sv"
`include "mem_mon.sv"
`include "mem_sqr.sv"
`include "mem_drv.sv"
`include "mem_agent.sv"
`include "mem_sbd.sv"
`include "mem_env.sv"
`include "seq_lib.sv"
`include "test_lib.sv"
`include "top.sv"

