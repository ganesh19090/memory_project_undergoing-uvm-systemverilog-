typedef uvm_sequencer#(mem_tx) mem_sqr;
//class mem_sqr extends uvm_sequencer;
////factory registration
//`uvm_component_utils(mem_sqr)
//
////new constructor
//function new (string name="",uvm_component parent);
//super.new(name,parent);
//endfunction
//
////build_phase
//function void build_phase(uvm_phase phase);
//$display("build_phase of mem_sqr is verified");
//endfunction
//
//endclass
