module top;
initial begin
run_test("mem_wr_rd_test");
end
endmodule
