module top;
initial begin
run_test("axi_test");
end
endmodule
