`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "mem_tx.sv"
`include "mem_wr_rd_seq.sv"
`include "mem_mon.sv"
`include "mem_sqr.sv"
`include "mem_drv.sv"
`include "mem_agent.sv"
`include "mem_env.sv"
`include "mem_wr_rd_test.sv"
`include "top.sv"

